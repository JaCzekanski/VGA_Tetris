��  CCircuit��  CSerializeHack           ��  CPart    h  h    ���  CEarth�� 	 CTerminal  ����       	                     ����         ��      �� 	 CVoltRail��  CValue  )37    5V(          @      �? V 
�  <0Q1              @�,�M�ɂ�    4,<4         ����     �
�  DHYI                            <:DR        ��      ��  CSPDT��  CToggle  hP�p        
�  �@�A              @�,�M�ɂ�  
�  X8m9              @�,�M�ɂ?  
�  XHmI      	                     l4�L         ��    �� 
 CVoltmeter��  CMeter  �Y�g      688(    
�  �@�U       	 K`�~��?          
�  �l��                            �T�l        ��      �
�  @-A      	         �,�M�ɂ?    ,44L    !    ��      �� 	 CResistor�  �.�<    470        `}@      �?   
�  �@�A        K`�~��?�,�M�ɂ�  
�  �@�A      	       @�,�M�ɂ?    �<�D    %    ��      "��  �.<    75        �R@      �?   
�  @A                �,�M�ɂ�  
�  �@�A      	 K`�~��?�,�M�ɂ?    �<D    )    ��      ��  CDiode
�  X�m�              @`zrV�xv?  
�  ����        )��b�T@`zrV�xv�    l���    -    ��      +�
�  X�m�              @`zrV�xv?  
�  ����        )��b�T@`zrV�xv�    l���    0    ��      +�
�  X�m�              @�ʺ[��s?  
�  ����        ���p�X@�ʺ[��s�    l���    3    ��      "��  ����    750        p�@      �?   
�  ����        A���?�ʺ[��s�  
�  ����      	 ���p�X@�ʺ[��s?    ����    7    ��      "��  ����    720        ��@      �?   
�  ����        W`r��?�zrV�xv�  
�  ����      	 )��b�T@�zrV�xv?    ����    ;    ��      "��  ����    720        ��@      �?   
�  ����        U`r��?�zrV�xv�  
�  ����      	 )��b�T@�zrV�xv?    ����    ?    ��      ��  0pP�     A   
�  L`aa              @��'Bs7��  
�   X5Y              @��'Bs7�?  
�   h5i                            4TLl    C     ��    �
�  h�}�     	                       |���    G    ��      ��  ,�T�      383   
�   �5�        W`r��?          
�  L�a�     	                       4�L    J   ��      ��  ,�T�      383   
�   �5�        U`r��?          
�  L�a�     	                       4�L�    N   ��      ��  ,�T�      688   
�   �5�        A���?          
�  L�a�     	                       4�L�    R   ��      ��  CVZero��  CText  � �     0V    
�  � �                 s/͹�I?    � �      X    ����     ��  � y� �    5V(          @      �? V 
�  � �� �              @��E�¡��    � |� �     [    ����     "��  ����    1k        @�@      �?k  
�  ����        W`r��?t/͹�9?  
�  ����      	         t/͹�9�    ����    ^    ��      "��  ����    1k        @�@      �?k  
�  ����        U`r��?r/͹�9?  
�  ����      	         r/͹�9�    ����    b    ��      "��  �F�T    1k        @�@      �?k  
�  �X�Y        A���?�"w$>�q�  
�  �X�Y     
 	       @�"w$>�q?    �T�\    f    ��      �
�  p���                !Ow�ٓ?    ����    i    ��      "��  (FHT    75        �R@      �?   
�  DXYY                ��@�ʂ�  
�  X-Y        A���?��@�ʂ?    ,TD\    l    ��      "��  (�H�    75        �R@      �?   
�  D�Y�                ���C�t�  
�  �-�        U`r��?���C�t?    ,�D�    p    ��      "��  (�H�    75        �R@      �?   
�  D�Y�                ���C�t�  
�  �-�        W`r��?���C�t?    ,�D�    t    ��      ��  p��      v   
�  ����                t/͹�9?  
�  `�u�              @          
�  `�u�                t/͹�9�    t���    x      ��    ��  p���      {   
�  ����                r/͹�9?  
�  `�u�              @          
�  `�u�                r/͹�9�    t���    }      ��    ��  ph��     �   
�  �X�Y     
         @�"w$>�q�  
�  `PuQ              @�"w$>�q?  
�  ``ua                            tL�d    �     ��        h  h    ���  CWire  X0Y9       ��  P0Y1      ��  X�Y�       ��  X�Y�       ��  X�Y�       ��  X�i�      ��  h`i�       ��  ``ia      ���� 
 CCrossOver  ����      ��  �T�\        ����       ����  ����      ��  �T�\        ����       ����  ����      ��  ����        ���Y       ����  ����      ��  ����        ����      ��  ����       ����  ����        ����      ��  ��!�      ��  ����       ��  ����      ��  � 8Q9      ��  � 8� 9      ����  � L� T        � h� 9       ��  � h!i      ����  � L� T        � PIQ      ��  � X� Q       ��  � X!Y      ����  N�T�        P`Q�       ��  P`aa      ��  HPaQ      ��  ���      ����  ����        ���      ����  �T�\      ��  �T�\        �XY      ��  ����      ��  ��!�      ��  ����      ��  ��!�      ��  `�a�      	 ��  `�a�      	 ��  `�i�     	 ��  `�a�      	 ��  � P� �       ��  � � 9       ��  P�Q9       ��  P�a�      ����  N�T�        P�Q�       ����  N�T�        H�a�      ��  P�a�      ����  N�T�        H�a�      ��  H�I�       ��  HPI�       ��  X�Y�       ��  X�Y�       ��  X�q�      ��  XXY�           h  h    �    h  h        h  h         �      &  �      %     ! ) ! % % * &  & ) ) ! *  * - � - . . < 0 � 0 1 1 @ 3 � 3 4 4 8 7 7 � 8 4 8 ; ; � < . < ? ? � @ 1 @ C C � D � D E � E G � G J � J K K � N � N O O � R � R S S � X X � [ [ � ^ ^ � _ x _ b b � c } c f f � g � g i � i l l � m � m p p � q � q t t � u � u x x _ y � y z � z } } c ~ � ~  �  � � g � � � � � � �   � 0 - 3 � � � � � � � C � � � � � � � � � � � � � � � � � � � � � � � ; � � � � � ? � � N � � 7 � � � � � � � � � � E � � � � � � � D � � � � � � � � � u � � � q � � � � f m ^ � � J b � � R � K O � � G S � � [ X � � � � z � � � � � � � y �  � � � ~ � � � � � t p � � i l �            �$s�        @     +        @            @    "V  (      ��                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 